//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 07/01/2023 09:54:34 PM
// Design Name: 
// Module Name: program_counter_add.sv
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module program_counter_add #(
  parameter DWIDTH = 32
)(
  input  logic [DWIDTH-1:0] Program_Count_Curr,	// Current Program Count
  output logic [DWIDTH-1:0] Program_Count_Next	  // Next Program Count
);

////////////////////////////////////////////////////////////////
///////////////////////   Module Logic   ///////////////////////
////////////////////////////////////////////////////////////////

always_comb begin
  Program_Count_Next <= Program_Count_Curr + 4;
end

////////////////////////////////////////////////////////////////
//////////////////   Instantiation Template   //////////////////
////////////////////////////////////////////////////////////////

/*
program_counter_add #(
  .DWIDTH()
)
program_counter_add (
  .Program_Count_Curr(),
  .Program_Count_Next()
);
*/

endmodule